// *****************************************************
// AVR address constants (localparams)
//  for registers used by Xcelerator Blocks (XBs) 
// *****************************************************

localparam LFSR_CTRL_Address = 8'he0;
localparam LFSR_SEED_Address = 8'he1;
localparam LFSR_DATA_Address = 8'he2;

